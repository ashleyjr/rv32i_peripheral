module x_top_mem#(
   p_clk_hz = 1000000, 
   p_baud   = 9600
)(
   input    logic          i_clk,
   input    logic          i_nrst,
   // Mem Interface
   input    logic          i_rnw,
   input    logic          i_valid,
   output   logic          o_accept,
   input    logic [31:0]   i_addr,
   input    logic [31:0]   i_data, 
   output   logic [31:0]   o_data,
   // UART Interface
   input    logic          i_rx,
   output   logic          o_tx
);

   typedef enum logic [6:0] {
      IDLE, 
      W_CMD,
      R_CMD,
      W0,
      R0, 
      W1,
      R1, 
      W2,
      R2, 
      W3,
      R3, 
      WD0,
      WD1,
      WD2,
      WD3,
      RD0,
      RD1,
      RD2,
      RD3
   } sm_t;
  
   logic    [7:0] tx_data; 
   logic          tx_valid;
   logic          tx_accept;

   logic    [7:0] rx_data;
   logic          rx_valid;
  
   sm_t           sm_d;
   sm_t           sm_q;
   logic          sm_en;

   logic          tx_valid_q;
   logic          tx_valid_d;

   logic          rx_ack;
   logic          rx_ack_d;
   logic          rx_ack_q;

   ///////////////////////////////////////////////////////////////////
   // State Machine

   assign sm_en = (sm_q == IDLE              ) ? i_valid: 
                  (sm_q inside {R_CMD, W_CMD}) ? tx_accept:
                                                 rx_ack;
                  
   always_comb begin
      case(sm_q) 
         IDLE:       if(i_rnw)   sm_d = R_CMD;
                     else        sm_d = W_CMD;
         R_CMD:                  sm_d = R0;
         R0:                     sm_d = R1; 
         R1:                     sm_d = R2; 
         R2:                     sm_d = R3; 
         R3:                     sm_d = RD0; 
         RD0:                    sm_d = RD0;
         RD1:                    sm_d = RD0;
         RD2:                    sm_d = RD0;
         RD3:                    sm_d = IDLE;
         W_CMD:                  sm_d = W0;
         W0:                     sm_d = W1; 
         W1:                     sm_d = W2; 
         W2:                     sm_d = W3; 
         W3:                     sm_d = WD0; 
         WD0:                    sm_d = WD0;
         WD1:                    sm_d = WD0;
         WD2:                    sm_d = WD0;
         WD3:                    sm_d = IDLE;
         default:                sm_d = IDLE;
      endcase
   end 

   always_ff@(posedge i_clk or negedge i_nrst) begin
      if(!i_nrst)    sm_q <= IDLE;
      else if(sm_en) sm_q <= sm_d;
   end 
   
   ///////////////////////////////////////////////////////////////////
   // Tx

   always_comb begin
      case(sm_q) 
         W_CMD:   tx_data = 8'b00000000;
         R_CMD:   tx_data = 8'h00000001; 
         W0,R0:   tx_data = i_addr[7:0];
         W1,R1:   tx_data = i_addr[15:8];
         W2,R2:   tx_data = i_addr[23:16];
         W3,R3:   tx_data = i_addr[31:24];
         WD0:     tx_data = i_data[7:0]; 
         WD1:     tx_data = i_data[15:8]; 
         WD2:     tx_data = i_data[23:16]; 
         WD3:     tx_data = i_data[31:24];
         default: tx_data = 'd0;
      endcase
   end

   assign tx_valid_d = sm_en | (tx_valid_q & ~tx_accept);

   always_ff@(posedge i_clk or negedge i_nrst) begin
      if(!i_nrst)    tx_valid_q <= 1'b0;
      else           tx_valid_q <= tx_valid_d;
   end 
   
   x_top_uart_tx #(
      .p_clk_hz   (p_clk_hz   ),
      .p_baud     (p_baud     )
   ) u_tx (
      .i_clk      (i_clk      ),
      .i_nrst     (i_nrst     ),
      .i_data     (tx_data    ),
      .o_tx       (o_tx       ),
      .i_valid    (tx_valid_q ),
      .o_accept   (tx_accept  )
   );

   ///////////////////////////////////////////////////////////////////
   // Rx

   assign rx_ack   = (rx_data == 'd0 & rx_valid); 
   assign rx_ack_d = (rx_ack_q) ? ~sm_en : rx_ack;   

   always_ff@(posedge i_clk or negedge i_nrst) begin
      if(!i_nrst)    rx_ack_q <= 1'b0;
      else           rx_ack_q <= rx_ack_d;
   end 
   
   x_top_uart_rx #(
      .p_clk_hz   (p_clk_hz   ),
      .p_baud     (p_baud     )
   ) u_rx (
      .i_clk      (i_clk      ),
      .i_nrst     (i_nrst     ),
      .i_rx       (i_rx       ),
      .o_valid    (rx_valid   ),
      .o_data     (rx_data    )
   );

endmodule
